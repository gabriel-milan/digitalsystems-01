----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:11:10 09/21/2018 
-- Design Name: 
-- Module Name:    XOR_4BITS - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity XOR_4BITS is
    Port ( A : in  STD_LOGIC_VECTOR(3 downto 0);
           --B : in  STD_LOGIC_VECTOR (3 downto 0);
           Z : out  STD_LOGIC_VECTOR(3 downto 0));
end XOR_4BITS;

architecture Behavioral of XOR_4BITS is

signal B : STD_LOGIC_VECTOR (3 downto 0);

begin
	
	B <= "1010";

	Z <= A xor B;
	
end Behavioral;

